module Decoder();

    
endmodule //moduleName


    


